
`timescale 1ps/1ps


module testbench;

    SYSC_FPGA
    i0_SYSC_FPGA
    (

	);

endmodule
