
`timescale 1ns/1ns


module testbench;

    SYSC_FPGA
    i0_SYSC_FPGA
    (

	);

endmodule
